--32-bit CPU