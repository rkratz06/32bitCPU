--alu controller